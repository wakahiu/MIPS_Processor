module ISR(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h27bdffec;
30'h00000001: inst = 32'hafbf0010;
30'h00000002: inst = 32'h401a6800;
30'h00000003: inst = 32'h401b6000;
30'h00000004: inst = 32'h00000000;
30'h00000005: inst = 32'h337bfc00;
30'h00000006: inst = 32'h035bd024;
30'h00000007: inst = 32'h335b8000;
30'h00000008: inst = 32'h1f60000a;
30'h00000009: inst = 32'h00000000;
30'h0000000a: inst = 32'h335b4000;
30'h0000000b: inst = 32'h1f60007d;
30'h0000000c: inst = 32'h00000000;
30'h0000000d: inst = 32'h335b0800;
30'h0000000e: inst = 32'h1f600086;
30'h0000000f: inst = 32'h00000000;
30'h00000010: inst = 32'h335b0400;
30'h00000011: inst = 32'h1f6000a3;
30'h00000012: inst = 32'h00000000;
30'h00000013: inst = 32'h3c1b1fff;
30'h00000014: inst = 32'h8f7a002c;
30'h00000015: inst = 32'h241b003c;
30'h00000016: inst = 32'h0c0000e2;
30'h00000017: inst = 32'h275a0001;
30'h00000018: inst = 32'h3c1b1fff;
30'h00000019: inst = 32'h8f7b0028;
30'h0000001a: inst = 32'h00000000;
30'h0000001b: inst = 32'h037ad021;
30'h0000001c: inst = 32'h3c1b1fff;
30'h0000001d: inst = 32'haf7a0028;
30'h0000001e: inst = 32'h8f7a002c;
30'h0000001f: inst = 32'h241b003c;
30'h00000020: inst = 32'h0c000103;
30'h00000021: inst = 32'h275a0001;
30'h00000022: inst = 32'h3c1b1fff;
30'h00000023: inst = 32'haf7a002c;
30'h00000024: inst = 32'h8f7a0024;
30'h00000025: inst = 32'h00000000;
30'h00000026: inst = 32'h1b400005;
30'h00000027: inst = 32'h00000000;
30'h00000028: inst = 32'h8f7a002c;
30'h00000029: inst = 32'h8f7b0028;
30'h0000002a: inst = 32'h0c000039;
30'h0000002b: inst = 32'h00000000;
30'h0000002c: inst = 32'h401b5800;
30'h0000002d: inst = 32'h3c1a02fa;
30'h0000002e: inst = 32'h375af080;
30'h0000002f: inst = 32'h035bd821;
30'h00000030: inst = 32'h409b5800;
30'h00000031: inst = 32'h00000000;
30'h00000032: inst = 32'h401b6800;
30'h00000033: inst = 32'h3c1affff;
30'h00000034: inst = 32'h375a7fff;
30'h00000035: inst = 32'h037ad824;
30'h00000036: inst = 32'h409b6800;
30'h00000037: inst = 32'h08000111;
30'h00000038: inst = 32'h00000000;
30'h00000039: inst = 32'h27bdffec;
30'h0000003a: inst = 32'hafa80010;
30'h0000003b: inst = 32'hafbf000c;
30'h0000003c: inst = 32'hafa90008;
30'h0000003d: inst = 32'h03404021;
30'h0000003e: inst = 32'h03604821;
30'h0000003f: inst = 32'h001bd021;
30'h00000040: inst = 32'h0c0000e2;
30'h00000041: inst = 32'h241b000a;
30'h00000042: inst = 32'h0c00005f;
30'h00000043: inst = 32'h275a0030;
30'h00000044: inst = 32'h241b000a;
30'h00000045: inst = 32'h0c000103;
30'h00000046: inst = 32'h0009d021;
30'h00000047: inst = 32'h0c00005f;
30'h00000048: inst = 32'h275a0030;
30'h00000049: inst = 32'h0c00005f;
30'h0000004a: inst = 32'h241a003a;
30'h0000004b: inst = 32'h0100d021;
30'h0000004c: inst = 32'h0c0000e2;
30'h0000004d: inst = 32'h241b000a;
30'h0000004e: inst = 32'h0c00005f;
30'h0000004f: inst = 32'h275a0030;
30'h00000050: inst = 32'h241b000a;
30'h00000051: inst = 32'h0c000103;
30'h00000052: inst = 32'h0008d021;
30'h00000053: inst = 32'h0c00005f;
30'h00000054: inst = 32'h275a0030;
30'h00000055: inst = 32'h0c00005f;
30'h00000056: inst = 32'h241a000d;
30'h00000057: inst = 32'h0c00005f;
30'h00000058: inst = 32'h241a000a;
30'h00000059: inst = 32'h8fa80010;
30'h0000005a: inst = 32'h8fa90008;
30'h0000005b: inst = 32'h8fbf000c;
30'h0000005c: inst = 32'h27bd0014;
30'h0000005d: inst = 32'h03e00008;
30'h0000005e: inst = 32'h00000000;
30'h0000005f: inst = 32'h27bdffe8;
30'h00000060: inst = 32'hafaa0014;
30'h00000061: inst = 32'hafbf0010;
30'h00000062: inst = 32'hafa8000c;
30'h00000063: inst = 32'hafa90008;
30'h00000064: inst = 32'hafba0004;
30'h00000065: inst = 32'hafbb0000;
30'h00000066: inst = 32'h3c1b8000;
30'h00000067: inst = 32'h8f7b0000;
30'h00000068: inst = 32'h00000000;
30'h00000069: inst = 32'h1f600015;
30'h0000006a: inst = 32'h00000000;
30'h0000006b: inst = 32'h3c081fff;
30'h0000006c: inst = 32'h8d1a0004;
30'h0000006d: inst = 32'h00000000;
30'h0000006e: inst = 32'h275a0001;
30'h0000006f: inst = 32'h0c000103;
30'h00000070: inst = 32'h241b0014;
30'h00000071: inst = 32'h8d090008;
30'h00000072: inst = 32'h03405021;
30'h00000073: inst = 32'h113a000d;
30'h00000074: inst = 32'h00000000;
30'h00000075: inst = 32'h8d1a0004;
30'h00000076: inst = 32'h2508000c;
30'h00000077: inst = 32'h0348d821;
30'h00000078: inst = 32'h8fa90004;
30'h00000079: inst = 32'h00000000;
30'h0000007a: inst = 32'ha3690000;
30'h0000007b: inst = 32'h0140d021;
30'h0000007c: inst = 32'h3c081fff;
30'h0000007d: inst = 32'h08000081;
30'h0000007e: inst = 32'had1a0004;
30'h0000007f: inst = 32'h3c1b8000;
30'h00000080: inst = 32'haf7a0008;
30'h00000081: inst = 32'h8faa0014;
30'h00000082: inst = 32'h8fbf0010;
30'h00000083: inst = 32'h8fa8000c;
30'h00000084: inst = 32'h8fa90008;
30'h00000085: inst = 32'h8fba0004;
30'h00000086: inst = 32'h8fbb0000;
30'h00000087: inst = 32'h03e00008;
30'h00000088: inst = 32'h27bd0018;
30'h00000089: inst = 32'h3c1b1fff;
30'h0000008a: inst = 32'h8f7a0000;
30'h0000008b: inst = 32'h00000000;
30'h0000008c: inst = 32'h275a0001;
30'h0000008d: inst = 32'haf7a0000;
30'h0000008e: inst = 32'h401b6800;
30'h0000008f: inst = 32'h3c1affff;
30'h00000090: inst = 32'h375abfff;
30'h00000091: inst = 32'h037ad824;
30'h00000092: inst = 32'h409b6800;
30'h00000093: inst = 32'h08000111;
30'h00000094: inst = 32'h00000000;
30'h00000095: inst = 32'h3c1a1fff;
30'h00000096: inst = 32'h8f5b0004;
30'h00000097: inst = 32'h8f5a0008;
30'h00000098: inst = 32'h00000000;
30'h00000099: inst = 32'h135b0014;
30'h0000009a: inst = 32'h00000000;
30'h0000009b: inst = 32'h3c1b1fff;
30'h0000009c: inst = 32'h277b000c;
30'h0000009d: inst = 32'h037ad821;
30'h0000009e: inst = 32'h837b0000;
30'h0000009f: inst = 32'h3c1a8000;
30'h000000a0: inst = 32'h8f5a0000;
30'h000000a1: inst = 32'h00000000;
30'h000000a2: inst = 32'h1b40000b;
30'h000000a3: inst = 32'h00000000;
30'h000000a4: inst = 32'h3c1a8000;
30'h000000a5: inst = 32'haf5b0008;
30'h000000a6: inst = 32'h3c1a1fff;
30'h000000a7: inst = 32'h8f5a0008;
30'h000000a8: inst = 32'h00000000;
30'h000000a9: inst = 32'h275a0001;
30'h000000aa: inst = 32'h0c000103;
30'h000000ab: inst = 32'h241b0014;
30'h000000ac: inst = 32'h3c1b1fff;
30'h000000ad: inst = 32'haf7a0008;
30'h000000ae: inst = 32'h401b6800;
30'h000000af: inst = 32'h3c1affff;
30'h000000b0: inst = 32'h375af7ff;
30'h000000b1: inst = 32'h037ad824;
30'h000000b2: inst = 32'h409b6800;
30'h000000b3: inst = 32'h08000111;
30'h000000b4: inst = 32'h00000000;
30'h000000b5: inst = 32'h3c1a8000;
30'h000000b6: inst = 32'h8f5b0004;
30'h000000b7: inst = 32'h00000000;
30'h000000b8: inst = 32'h1b600058;
30'h000000b9: inst = 32'h00000000;
30'h000000ba: inst = 32'h8f5a000c;
30'h000000bb: inst = 32'h0c00005f;
30'h000000bc: inst = 32'h00000000;
30'h000000bd: inst = 32'h241b0065;
30'h000000be: inst = 32'h137a0012;
30'h000000bf: inst = 32'h00000000;
30'h000000c0: inst = 32'h241b0064;
30'h000000c1: inst = 32'h137a0013;
30'h000000c2: inst = 32'h00000000;
30'h000000c3: inst = 32'h241b0072;
30'h000000c4: inst = 32'h137a0013;
30'h000000c5: inst = 32'h00000000;
30'h000000c6: inst = 32'h241b0052;
30'h000000c7: inst = 32'h137a0010;
30'h000000c8: inst = 32'h00000000;
30'h000000c9: inst = 32'h241b0076;
30'h000000ca: inst = 32'h137a000d;
30'h000000cb: inst = 32'h00000000;
30'h000000cc: inst = 32'h241b0056;
30'h000000cd: inst = 32'h137a000a;
30'h000000ce: inst = 32'h00000000;
30'h000000cf: inst = 32'h080000db;
30'h000000d0: inst = 32'h00000000;
30'h000000d1: inst = 32'h3c1b1fff;
30'h000000d2: inst = 32'h241a0001;
30'h000000d3: inst = 32'h080000db;
30'h000000d4: inst = 32'haf7a0024;
30'h000000d5: inst = 32'h3c1b1fff;
30'h000000d6: inst = 32'h080000db;
30'h000000d7: inst = 32'haf600024;
30'h000000d8: inst = 32'h3c1a1fff;
30'h000000d9: inst = 32'h080000db;
30'h000000da: inst = 32'haf5b0020;
30'h000000db: inst = 32'h401b6800;
30'h000000dc: inst = 32'h3c1affff;
30'h000000dd: inst = 32'h375afbff;
30'h000000de: inst = 32'h037ad824;
30'h000000df: inst = 32'h409b6800;
30'h000000e0: inst = 32'h08000111;
30'h000000e1: inst = 32'h00000000;
30'h000000e2: inst = 32'h27bdffec;
30'h000000e3: inst = 32'hafbf0010;
30'h000000e4: inst = 32'hafa4000c;
30'h000000e5: inst = 32'hafa80008;
30'h000000e6: inst = 32'h00002024;
30'h000000e7: inst = 32'h035b402b;
30'h000000e8: inst = 32'h1d000004;
30'h000000e9: inst = 32'h00000000;
30'h000000ea: inst = 32'h035bd023;
30'h000000eb: inst = 32'h080000e7;
30'h000000ec: inst = 32'h24840001;
30'h000000ed: inst = 32'h0080d021;
30'h000000ee: inst = 32'h8fbf0010;
30'h000000ef: inst = 32'h8fa4000c;
30'h000000f0: inst = 32'h8fa80008;
30'h000000f1: inst = 32'h03e00008;
30'h000000f2: inst = 32'h27bd0014;
30'h000000f3: inst = 32'h27bdffec;
30'h000000f4: inst = 32'hafbf0010;
30'h000000f5: inst = 32'hafa4000c;
30'h000000f6: inst = 32'hafa80008;
30'h000000f7: inst = 32'h00002024;
30'h000000f8: inst = 32'h13600004;
30'h000000f9: inst = 32'h00000000;
30'h000000fa: inst = 32'h277bffff;
30'h000000fb: inst = 32'h080000f8;
30'h000000fc: inst = 32'h009a2021;
30'h000000fd: inst = 32'h0080d021;
30'h000000fe: inst = 32'h8fbf0010;
30'h000000ff: inst = 32'h8fa4000c;
30'h00000100: inst = 32'h8fa80008;
30'h00000101: inst = 32'h03e00008;
30'h00000102: inst = 32'h27bd0014;
30'h00000103: inst = 32'h27bdffec;
30'h00000104: inst = 32'hafbf0010;
30'h00000105: inst = 32'hafa4000c;
30'h00000106: inst = 32'hafa80008;
30'h00000107: inst = 32'h035b402b;
30'h00000108: inst = 32'h1d000003;
30'h00000109: inst = 32'h00000000;
30'h0000010a: inst = 32'h08000107;
30'h0000010b: inst = 32'h035bd023;
30'h0000010c: inst = 32'h8fbf0010;
30'h0000010d: inst = 32'h8fa4000c;
30'h0000010e: inst = 32'h8fa80008;
30'h0000010f: inst = 32'h03e00008;
30'h00000110: inst = 32'h27bd0014;
30'h00000111: inst = 32'h8fbf0010;
30'h00000112: inst = 32'h27bd0014;
30'h00000113: inst = 32'h401a7000;
30'h00000114: inst = 32'h401b6000;
30'h00000115: inst = 32'h00000000;
30'h00000116: inst = 32'h377b0001;
30'h00000117: inst = 32'h409b6000;
30'h00000118: inst = 32'h03400008;
30'h00000119: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
