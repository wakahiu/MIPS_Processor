module game(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c000003;
30'h00000002: inst = 32'h37bd1000;
30'h00000003: inst = 32'h27bdffe8;
30'h00000004: inst = 32'h3c028000;
30'h00000005: inst = 32'h3c031040;
30'h00000006: inst = 32'h3c0410c0;
30'h00000007: inst = 32'h34450010;
30'h00000008: inst = 32'h34630000;
30'h00000009: inst = 32'hafa00010;
30'h0000000a: inst = 32'h3c060100;
30'h0000000b: inst = 32'h34870000;
30'h0000000c: inst = 32'h34480014;
30'h0000000d: inst = 32'haca30000;
30'h0000000e: inst = 32'h3c0302ff;
30'h0000000f: inst = 32'h34c600ff;
30'h00000010: inst = 32'had070000;
30'h00000011: inst = 32'h3c08000a;
30'h00000012: inst = 32'h34630000;
30'h00000013: inst = 32'h34890004;
30'h00000014: inst = 32'hace60000;
30'h00000015: inst = 32'h3c060315;
30'h00000016: inst = 32'h3507000a;
30'h00000017: inst = 32'h34880008;
30'h00000018: inst = 32'had230000;
30'h00000019: inst = 32'h34c3000a;
30'h0000001a: inst = 32'h3486000c;
30'h0000001b: inst = 32'had070000;
30'h0000001c: inst = 32'h3c071080;
30'h0000001d: inst = 32'h34840010;
30'h0000001e: inst = 32'hacc30000;
30'h0000001f: inst = 32'h34e30000;
30'h00000020: inst = 32'h34460018;
30'h00000021: inst = 32'hac800000;
30'h00000022: inst = 32'h24040001;
30'h00000023: inst = 32'h3442001c;
30'h00000024: inst = 32'hacc30000;
30'h00000025: inst = 32'hac440000;
30'h00000026: inst = 32'haca30000;
30'h00000027: inst = 32'h8fa20010;
30'h00000028: inst = 32'h00000000;
30'h00000029: inst = 32'h27bd0018;
30'h0000002a: inst = 32'h03e00008;
30'h0000002b: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
